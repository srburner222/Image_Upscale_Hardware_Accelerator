 localparam HRES = 128;
 localparam VRES = 128;