/**
 * BSG Test Node Client
 */

/**********
 * NOTICE *
 **********
 * This file has been modified from its original form found in:
 * https://github.com/bsg-external/ee478-designs-project
 * 
 * This file is subject to the license found at the following link:
 * http://solderpad.org/licenses/SHL-0.51
 * 
 * Further licensing details can be found in the repo linked above
 */

module  bsg_test_node_client #(parameter ring_width_p="inv"
                              ,parameter master_p="inv"
                              ,parameter master_id_p="inv"
                              ,parameter client_id_p="inv")
  (input  clk_i
  ,input  reset_i
  ,input  en_i

  ,input                     v_i
  ,input  [ring_width_p-1:0] data_i
  ,output                    ready_o
  
  ,output                    v_o
  ,output [ring_width_p-1:0] data_o
  ,input                     yumi_i
  );

   // Include image scale parameters generated by runsim.py
  `include "v/parameters.vh"
   
  logic [74:0] data_li;
  logic [31:0] data_lo;
   
  assign data_li = data_i[74:0];
  assign data_o  = { 4'(client_id_p), {51{1'b0}}, data_lo };

  /** INSTANTIATE NODE 0 **/
  if ( client_id_p == 0 ) begin

     interpolation #(.bit_depth(8), .v_res(VRES), .h_res(HRES)) 
                   interpolate_r (.clk       (clk_i),
			          .reset     (reset_i),
				  .valid_in  (v_i),
				  .data_in   (data_li[23:16]),
				  .valid_out (v_o),
				  .ready_out (ready_o),
				  .data_out  (data_lo[23:16])
				 );

     interpolation #(.bit_depth(8), .v_res(VRES), .h_res(HRES)) 
                   interpolate_g (.clk       (clk_i),
			          .reset     (reset_i),
				  .valid_in  (v_i),
				  .data_in   (data_li[15:8]),
				  .valid_out (v_o),
				  .ready_out (ready_o),
				  .data_out  (data_lo[15:8])
				 );

     interpolation #(.bit_depth(8), .v_res(VRES), .h_res(HRES)) 
                   interpolate_b (.clk       (clk_i),
			          .reset     (reset_i),
				  .valid_in  (v_i),
				  .data_in   (data_li[7:0]),
				  .valid_out (v_o),
				  .ready_out (ready_o),
				  .data_out  (data_lo[7:0])
				 );
     
  end
  /** INSTANTIATE NODE 1 **/
//  else if ( client_id_p == 1 ) begin
//
//    <INSTANTIATE NODE MODULE>
//
//  end

endmodule

